`default_nettype none
`timescale 1ns/1ns
module debounce
(
    input wire clk,
    input wire reset,
    input wire button,
    output reg debounced
);

endmodule
