`default_nettype none
`timescale 1ns/1ns
module rgb_mixer (
    input clk,
    input reset_n,
    input enc0_a,
    input enc0_b,
    input enc1_a,
    input enc1_b,
    input enc2_a,
    input enc2_b,
    output pwm0_out,
    output pwm1_out,
    output pwm2_out
);

endmodule
