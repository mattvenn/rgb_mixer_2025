`default_nettype none
`timescale 1ns/1ns
module pwm (
    input wire clk,
    input wire reset,
    output reg out,
    input wire [7:0] level
    );

endmodule
